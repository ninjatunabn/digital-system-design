library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Johnson_Counter is
    Port (Clock, Reset : in  STD_LOGIC;
        Q     : out STD_LOGIC_VECTOR(7 downto 0));
end Johnson_Counter;

architecture Behavioral of Johnson_Counter is
    signal count : STD_LOGIC_VECTOR(7 downto 0) := "00000000";
begin
    process(Clock, Reset)
    begin
        if Reset = '1' then
            count <= "00000000";
        elsif rising_edge(Clock) then
            count <= count(6 downto 0) & not count(7);
        end if;
    end process;
    Q <= count;
end Behavioral;
